// 853355 Davi Puddo

// constant definitions
`define found 1
`define notfound 0

// Definir clock
module clock (clk);

	output reg clk;

	initial
		begin
			clk = 1'b0;
		end
	
	always
		begin
			#1 clk = ~clk;
		end

endmodule // clock

// FSM by Mealy
module mealy ( y, x, clk, reset );

	output y;
	input x;
	input clk;
	input reset;
	reg y;

	parameter // state identifiers
	start = 2'b00,
	id1 = 2'b01,
	id11 = 2'b11,
	id110 = 2'b10;
	reg [1:0] E1; // current state variables
	reg [1:0] E2; // next state logic output
	// next state logic
	always @( x or E1 )
	begin
		y = `notfound;
		case ( E1 )
			start:
				if ( x )
					E2 = id1;
				else
					E2 = start;
			id1:
				if ( x )
					E2 = id11;
				else
					E2 = start;
			id11:
				if ( x )
					E2 = id11;
				else
					E2 = id110;
			id110:
				if ( x )
					begin
						E2 = id1;
						y = `found;
					end
				else
					begin
						E2 = start;
						y = `notfound;
					end
			default: // undefined state
				E2 = 2'bxx;
		endcase
	end // always at signal or state changing

	// state variables
	always @( posedge clk or negedge reset )
	begin
		if ( reset )
			E1 = E2; // updates current state
		else
			E1 = 0; // reset
	end // always at signal changing

endmodule // mealy

module G1101;

	// Definir dados
	reg x = 1'b0;
	reg reset = 1'b0;
	wire clk;
	wire y;

	// Chamar modulos
	clock C1 (clk);
	mealy M1 (y, x, clk, reset);

	always @(clk)
		#2 $display ("x: %b", x);

		initial
			begin : main

				#2 x = 1'b0; reset = 1'b1;
				#2 x = 1'b1; // 1
				#2 x = 1'b1; // 1
				#2 x = 1'b0; // 0
				#2 x = 1'b1; // 1
				#2 x = 1'b0;
				#2 x = 1'b1;
				#2 x = 1'b1; // 1
				#2 x = 1'b1; // 1
				#2 x = 1'b0; // 0
				#2 x = 1'b1; // 1

				#0 $finish;
			end // main
	
	// Mostrar resultado
	always @(posedge y)
		$display ("encontrado");

endmodule // G1101
